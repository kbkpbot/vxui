module vxui

import time

// =============================================================================
// Error Type Tests
// =============================================================================

fn test_vxui_error_enum() {
	assert int(VxuiError.unknown) == 0
	assert int(VxuiError.client_not_found) == 1
	assert int(VxuiError.no_clients) == 2
	assert int(VxuiError.no_valid_connection) == 3
	assert int(VxuiError.js_timeout) == 4
	assert int(VxuiError.js_validation_failed) == 5
}

fn test_vxui_error_detail_struct() {
	err := VxuiErrorDetail{
		code:    VxuiError.client_not_found
		message: 'Client not found'
		details: {
			'client_id': 'test-123'
		}
	}
	assert err.code == VxuiError.client_not_found
	assert err.message == 'Client not found'
	assert err.details['client_id'] == 'test-123'
}

fn test_vxui_error_detail_str() {
	err := VxuiErrorDetail{
		code:    VxuiError.auth_failed
		message: 'Authentication failed'
	}
	assert err.str() == 'Authentication failed'
}

fn test_new_error_detail() {
	err := new_error_detail(VxuiError.no_clients, 'No connected clients')
	assert err.code == VxuiError.no_clients
	assert err.message == 'No connected clients'
}

fn test_new_error_detail_with_details() {
	err := new_error_detail_with_details(VxuiError.client_not_found, 'Client not found',
		{
		'id': 'abc'
	})
	assert err.code == VxuiError.client_not_found
	assert err.details['id'] == 'abc'
}

// =============================================================================
// Event System Tests
// =============================================================================

fn test_event_type_enum() {
	assert int(EventType.before_start) == 0
	assert int(EventType.after_start) == 1
	assert int(EventType.client_connecting) == 2
	assert int(EventType.client_connected) == 3
	assert int(EventType.client_disconnected) == 4
	assert int(EventType.before_shutdown) == 5
	assert int(EventType.error) == 6
	assert int(EventType.js_execution) == 7
	assert int(EventType.before_request) == 8
	assert int(EventType.after_request) == 9
	assert int(EventType.middleware_error) == 10
}

fn test_event_data_struct() {
	data := EventData{
		event_type: EventType.client_connected
		client_id:  'test-client'
		message:    'Client connected'
	}
	assert data.event_type == EventType.client_connected
	assert data.client_id == 'test-client'
}

// =============================================================================
// Request/Response Tests
// =============================================================================

fn test_verb_enum() {
	assert int(Verb.any_verb) == 0
	assert int(Verb.get) == 1
	assert int(Verb.post) == 2
	assert int(Verb.put) == 3
	assert int(Verb.delete) == 4
	assert int(Verb.patch) == 5
}

fn test_request_struct() {
	req := Request{
		id:         'req-123'
		verb:       Verb.post
		path:       '/api/test'
		parameters: {
			'key': 'value'
		}
		headers:    {
			'Content-Type': 'application/json'
		}
		body:       '{"test": true}'
		client_id:  'client-1'
	}
	assert req.id == 'req-123'
	assert req.verb == Verb.post
	assert req.path == '/api/test'
	assert req.parameters['key'] == 'value'
}

fn test_response_struct() {
	mut resp := Response{
		status: 200
		body:   '{"result": "ok"}'
	}
	assert resp.status == 200
	assert resp.body == '{"result": "ok"}'

	resp.status = 404
	assert resp.status == 404
}

fn test_response_default_status() {
	resp := Response{}
	assert resp.status == 200
}

// =============================================================================
// Middleware Tests
// =============================================================================

fn test_middleware_context_struct() {
	req := Request{
		id:   'req-1'
		verb: Verb.get
		path: '/test'
	}
	mctx := MiddlewareContext{
		request:  req
		response: Response{}
	}
	assert mctx.request.id == 'req-1'
	assert mctx.response.status == 200
}

fn test_middleware_result_enum() {
	assert int(MiddlewareResult.continue_) == 0
	assert int(MiddlewareResult.stop) == 1
	assert int(MiddlewareResult.error) == 2
}

// =============================================================================
// Configuration Tests
// =============================================================================

fn test_config_defaults() {
	config := Config{}
	assert config.close_timer_ms == 5000
	assert config.ws_ping_interval_ms == 30000
	assert config.ws_pong_timeout_ms == 60000
	assert config.require_auth == true
	assert config.multi_client == false
	assert config.max_clients == 10
	assert config.js_timeout == 5000
	assert config.js_poll_ms == 10
	assert config.app_name == 'vxui-app'
}

fn test_config_custom() {
	config := Config{
		app_name:       'my-app'
		close_timer_ms: 10000
		multi_client:   true
		max_clients:    5
		window:         WindowConfig{
			width:  1920
			height: 1080
		}
	}
	assert config.app_name == 'my-app'
	assert config.close_timer_ms == 10000
	assert config.multi_client == true
	assert config.max_clients == 5
	assert config.window.width == 1920
}

fn test_js_sandbox_config_defaults() {
	config := JsSandboxConfig{}
	assert config.enabled == true
	assert config.timeout_ms == 5000
	assert config.max_result_size == 1048576
	assert config.allow_eval == false
	assert config.allowed_apis.len > 0
	assert config.forbidden_patterns.len > 0
}

fn test_js_sandbox_config_custom() {
	config := JsSandboxConfig{
		enabled:         false
		timeout_ms:      10000
		max_result_size: 2097152
		allow_eval:      true
	}
	assert config.enabled == false
	assert config.timeout_ms == 10000
	assert config.max_result_size == 2097152
	assert config.allow_eval == true
}

fn test_window_config_defaults() {
	config := WindowConfig{}
	assert config.width == 800
	assert config.height == 600
	assert config.x == -1
	assert config.y == -1
	assert config.resizable == true
}

fn test_window_config_custom() {
	config := WindowConfig{
		width:     1920
		height:    1080
		x:         100
		y:         50
		resizable: false
		title:     'My App'
	}
	assert config.width == 1920
	assert config.height == 1080
	assert config.title == 'My App'
}

fn test_browser_config_defaults() {
	config := BrowserConfig{}
	assert config.custom_args.len == 0
	assert config.headless == false
	assert config.devtools == false
	assert config.no_sandbox == false
}

fn test_browser_config_custom() {
	config := BrowserConfig{
		custom_args: ['--test-arg']
		headless:    true
		devtools:    true
		no_sandbox:  true
	}
	assert config.custom_args.len == 1
	assert config.headless == true
	assert config.devtools == true
	assert config.no_sandbox == true
}

fn test_reconnect_config_defaults() {
	config := ReconnectConfig{}
	assert config.enabled == true
	assert config.max_attempts == 5
	assert config.base_delay_ms == 1000
	assert config.max_delay_ms == 30000
	assert config.strategy == BackoffStrategy.full_jitter
}

fn test_reconnect_config_custom() {
	config := ReconnectConfig{
		enabled:       false
		max_attempts:  10
		base_delay_ms: 2000
		strategy:      BackoffStrategy.exponential
	}
	assert config.enabled == false
	assert config.max_attempts == 10
	assert config.strategy == BackoffStrategy.exponential
}

fn test_rate_limit_config_defaults() {
	config := RateLimitConfig{}
	assert config.enabled == true
	assert config.max_requests == 100
	assert config.window_ms == 60000
	assert config.block_duration == 30000
}

fn test_rate_limit_config_custom() {
	config := RateLimitConfig{
		enabled:      false
		max_requests: 50
		window_ms:    30000
	}
	assert config.enabled == false
	assert config.max_requests == 50
	assert config.window_ms == 30000
}

fn test_request_config_defaults() {
	config := RequestConfig{}
	assert config.timeout_ms == 30000
	assert config.retry_count == 0
	assert config.retry_delay_ms == 1000
}

fn test_log_config_defaults() {
	config := LogConfig{}
	assert config.level == .info
	assert config.output == 'stderr'
	assert config.max_file_size == 10485760
	assert config.rotate_files == 5
}

// =============================================================================
// Client Tests
// =============================================================================

fn test_client_struct() {
	now := time.now()
	client := Client{
		id:            'test-client-123'
		token:         'secret-token'
		connected:     now
		last_ping:     now
		request_count: 5
	}
	assert client.id == 'test-client-123'
	assert client.token == 'secret-token'
	assert client.request_count == 5
	assert client.connection == none
}

// =============================================================================
// Context Tests
// =============================================================================

fn test_context_defaults() {
	ctx := Context{}
	assert ctx.close_timer_ms == 5000
	assert ctx.js_poll_ms == 10
	assert ctx.multi_client == false
	assert ctx.clients.len == 0
}

fn test_context_with_config() {
	mut ctx := Context{}
	ctx.config = Config{
		app_name:       'test-app'
		close_timer_ms: 8000
	}
	assert ctx.config.app_name == 'test-app'
	assert ctx.config.close_timer_ms == 8000
}

fn test_get_clients_empty() {
	mut ctx := Context{}
	clients := ctx.get_clients()
	assert clients.len == 0
}

fn test_get_client_count_empty() {
	mut ctx := Context{}
	count := ctx.get_client_count()
	assert count == 0
}

fn test_get_port_initial() {
	ctx := Context{}
	assert ctx.get_port() == 0
}

fn test_get_token_initial() {
	ctx := Context{}
	assert ctx.get_token() == ''
}

fn test_get_token_custom() {
	mut ctx := Context{}
	ctx.token = 'my-secret-token'
	assert ctx.get_token() == 'my-secret-token'
}

fn test_get_config() {
	mut ctx := Context{}
	ctx.config = Config{
		app_name: 'test'
	}
	config := ctx.get_config()
	assert config.app_name == 'test'
}

// =============================================================================
// Setter Tests
// =============================================================================

fn test_set_window_size() {
	mut ctx := Context{}
	ctx.set_window_size(1024, 768)
	assert ctx.window.width == 1024
	assert ctx.window.height == 768
}

fn test_set_window_position() {
	mut ctx := Context{}
	ctx.set_window_position(100, 200)
	assert ctx.window.x == 100
	assert ctx.window.y == 200
}

fn test_set_window_title() {
	mut ctx := Context{}
	ctx.set_window_title('My Application')
	assert ctx.window.title == 'My Application'
}

fn test_set_resizable() {
	mut ctx := Context{}
	ctx.set_resizable(false)
	assert ctx.window.resizable == false
}

fn test_set_js_sandbox() {
	mut ctx := Context{}
	config := JsSandboxConfig{
		timeout_ms: 3000
	}
	ctx.set_js_sandbox(config)
	assert ctx.js_sandbox.timeout_ms == 3000
}

fn test_set_browser_config() {
	mut ctx := Context{}
	config := BrowserConfig{
		headless: true
	}
	ctx.set_browser_config(config)
	assert ctx.browser.headless == true
}

fn test_set_rate_limit() {
	mut ctx := Context{}
	config := RateLimitConfig{
		max_requests: 50
	}
	ctx.set_rate_limit(config)
	assert ctx.config.rate_limit.max_requests == 50
}

// =============================================================================
// Client Management Error Tests
// =============================================================================

fn test_close_client_not_found() {
	mut ctx := Context{}
	ctx.close_client('non-existent-id') or {
		assert err.msg().contains('not found')
		return
	}
	assert false
}

fn test_send_to_client_not_found() {
	mut ctx := Context{}
	ctx.send_to_client('non-existent-id', 'test') or {
		assert err.msg().contains('not found')
		return
	}
	assert false
}

fn test_ping_client_not_found() {
	mut ctx := Context{}
	ctx.ping_client('non-existent-id') or {
		assert err.msg().contains('not found')
		return
	}
	assert false
}

fn test_run_js_no_clients() {
	mut ctx := Context{}
	ctx.run_js('alert(1)', 1000) or {
		assert err.msg().contains('No connected clients')
		return
	}
	assert false
}

fn test_run_js_client_not_found() {
	mut ctx := Context{}
	ctx.run_js_client('non-existent-id', 'alert(1)', 1000) or {
		assert err.msg().contains('No connected clients') || err.msg().contains('not found')
		return
	}
	assert false
}

fn test_get_client_not_found() {
	mut ctx := Context{}
	client := ctx.get_client('non-existent-id')
	assert client == none
}

// =============================================================================
// Broadcast Tests
// =============================================================================

fn test_broadcast_no_clients() {
	mut ctx := Context{}
	ctx.broadcast('test message') or { return }
}

fn test_broadcast_except_no_clients() {
	mut ctx := Context{}
	ctx.broadcast_except('test message', 'client-1') or { return }
}

fn test_ping_all_clients_no_clients() {
	mut ctx := Context{}
	ctx.ping_all_clients()
}

// =============================================================================
// JS Validation Tests
// =============================================================================

fn test_validate_js_code_safe() {
	sandbox := JsSandboxConfig{
		enabled:            true
		forbidden_patterns: ['eval(', 'fetch(']
	}

	validate_js_code('document.title', sandbox) or {
		assert false
		return
	}
}

fn test_validate_js_code_forbidden() {
	sandbox := JsSandboxConfig{
		enabled:            true
		forbidden_patterns: ['eval(', 'fetch(']
	}

	validate_js_code('eval("alert(1)")', sandbox) or {
		assert err.msg().contains('Forbidden pattern')
		return
	}
	assert false
}

// =============================================================================
// Verb Strings Map Tests
// =============================================================================

fn test_verb_strings_map() {
	assert 'get' in verb_strings
	assert 'post' in verb_strings
	assert 'put' in verb_strings
	assert 'delete' in verb_strings
	assert 'patch' in verb_strings

	assert verb_strings['get'] == Verb.get
	assert verb_strings['post'] == Verb.post
}

// =============================================================================
// Route Tests
// =============================================================================

fn test_route_struct() {
	route := Route{
		verb: [Verb.get, Verb.post]
		path: '/api/test'
	}
	assert route.path == '/api/test'
	assert route.verb.len == 2
	assert Verb.get in route.verb
}

fn test_parse_attrs_empty() {
	verbs, path := parse_attrs('test', []) or {
		assert false
		return
	}
	assert path == '/test'
	assert verbs.len == 1
	assert Verb.any_verb in verbs
}

fn test_parse_attrs_with_path() {
	verbs, path := parse_attrs('test', ['/custom']) or {
		assert false
		return
	}
	assert path == '/custom'
}

fn test_parse_attrs_with_verb() {
	verbs, path := parse_attrs('test', ['get', 'post']) or {
		assert false
		return
	}
	assert verbs.len == 2
	assert Verb.get in verbs
	assert Verb.post in verbs
}

fn test_parse_attrs_duplicate_path() {
	parse_attrs('test', ['/path1', '/path2']) or { return }
	assert false
}

fn test_parse_attrs_invalid_verb() {
	parse_attrs('test', ['invalid_verb']) or { return }
	assert false
}

// =============================================================================
// Utility Tests
// =============================================================================

fn test_get_free_port() {
	port := get_free_port() or {
		assert false
		return
	}
	assert port >= 1025 && port <= 65534
}

fn test_sanitize_path_valid() {
	valid_paths := ['./ui/index.html', 'static/page.html', 'file.txt']
	for path in valid_paths {
		sanitize_path(path) or {
			assert false
			return
		}
	}
}

fn test_sanitize_path_traversal() {
	invalid_paths := ['../etc/passwd', '~/secret.txt', '/absolute/path']
	for path in invalid_paths {
		sanitize_path(path) or { continue }
		assert false
	}
}

fn test_escape_html() {
	assert escape_html('<script>') == '&lt;script&gt;'
	assert escape_html('"quoted"') == '&quot;quoted&quot;'
	assert escape_html('a & b') == 'a &amp; b'
}

fn test_escape_js() {
	assert escape_js('"quoted"') == '\\"quoted\\"'
	assert escape_js('line\nbreak') == 'line\\nbreak'
}

fn test_escape_attr() {
	assert escape_attr('"value"') == '&quot;value&quot;'
	assert escape_attr('a & b') == 'a &amp; b'
}

fn test_truncate_string() {
	assert truncate_string('hello', 10) == 'hello'
	assert truncate_string('hello world', 8) == 'hello...'
}

fn test_is_valid_email() {
	assert is_valid_email('test@example.com') == true
	assert is_valid_email('invalid') == false
}

fn test_generate_id() {
	id1 := generate_id()
	id2 := generate_id()
	assert id1.len == 16
	assert id1 != id2
}

// =============================================================================
// PackedApp Tests
// =============================================================================

fn test_packed_app_new() {
	packed := new_packed_app()
	assert packed.files.len == 0
	assert packed.total_size() == 0
}

fn test_packed_app_add_file() {
	mut packed := new_packed_app()
	packed.add_file('test.html', 'Hello'.bytes())
	assert packed.files.len == 1
	assert packed.has_file('test.html')
	assert packed.total_size() == 5
}

fn test_packed_app_add_file_string() {
	mut packed := new_packed_app()
	packed.add_file_string('index.html', '<html></html>')
	assert packed.files.len == 1

	content := packed.get_file_content('index.html')!
	assert content == '<html></html>'
}

fn test_packed_app_get_file_not_found() {
	packed := new_packed_app()
	packed.get_file('nonexistent') or {
		assert err.msg().contains('not found')
		return
	}
	assert false
}

fn test_packed_app_list_files() {
	mut packed := new_packed_app()
	packed.add_file_string('a.html', 'a')
	packed.add_file_string('b.css', 'b')

	files := packed.list_files()
	assert files.len == 2
}

// =============================================================================
// BackoffStrategy Tests
// =============================================================================

fn test_backoff_strategy_enum() {
	assert int(BackoffStrategy.constant) == 0
	assert int(BackoffStrategy.linear) == 1
	assert int(BackoffStrategy.exponential) == 2
	assert int(BackoffStrategy.full_jitter) == 3
}

// =============================================================================
// on_event Test
// =============================================================================

fn test_on_event() {
	mut ctx := Context{}
	ctx.on_event(EventType.client_connected, fn (e EventData) {
		// Handler registered
	})
	assert ctx.event_handlers[EventType.client_connected].len == 1
}

// =============================================================================
// use Middleware Test
// =============================================================================

fn test_use_middleware() {
	mut ctx := Context{}
	ctx.use(fn (mut mctx MiddlewareContext) MiddlewareResult {
		return .continue_
	})
	assert ctx.middlewares.len == 1
}
